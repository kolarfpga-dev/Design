//Basic top module that can be used to get utilization estimates
//Instantiate modules inside of this 
module basic_top(
    input logic clk,
    input logic rst,
    input logic in,
    output logic out
);
endmodule