//Macros for the sra(Simple Register Access) Interface